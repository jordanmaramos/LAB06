library verilog;
use verilog.vl_types.all;
entity contadordec_vlg_vec_tst is
end contadordec_vlg_vec_tst;
